library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity generic_uart is
    generic (
    );
    port (
    );
end entity generic_uart;

architecture Behavioral of generic_uart is
end architecture Behavioral;

